module cpu(
        inout [7:0] main_bus,
        input rst,
        input clk,
        input iclk,

        output [3:0] fout,

        /* verilator lint_off UNUSED */
        input [31:0] control_word
    );

    /* verilator lint_off PINMISSING */
    cword_splitter splitter(.control_word(control_word));
    alu_block alu(.main_bus(main_bus), .rst(rst), .clk(clk), .iclk(iclk), .fout(fout),
        .outctl(splitter.outctl),
        .loadctl(splitter.loadctl),
        .arg_l(splitter.alu_arg_l),
        .arg_r(splitter.alu_arg_r),
        .alt(splitter.alu_alt),
        .calcfn(splitter.flags_calc),
        .cin(splitter.carry));

endmodule
